// The configuration file of the DUT

`define DUT_WIDTH 4
